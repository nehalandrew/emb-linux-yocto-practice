module tb()
{
    return 0;
}